magic
tech sky130A
timestamp 1712479693
<< nwell >>
rect 0 -50 275 420
<< nmos >>
rect 130 -200 145 -100
<< pmos >>
rect 130 -5 145 205
<< ndiff >>
rect 85 -110 130 -100
rect 85 -190 95 -110
rect 115 -190 130 -110
rect 85 -200 130 -190
rect 145 -110 190 -100
rect 145 -190 160 -110
rect 180 -190 190 -110
rect 145 -200 190 -190
<< pdiff >>
rect 80 195 130 205
rect 80 5 90 195
rect 115 5 130 195
rect 80 -5 130 5
rect 145 195 195 205
rect 145 5 160 195
rect 185 5 195 195
rect 145 -5 195 5
<< ndiffc >>
rect 95 -190 115 -110
rect 160 -190 180 -110
<< pdiffc >>
rect 90 5 115 195
rect 160 5 185 195
<< psubdiff >>
rect 80 -250 195 -235
rect 80 -280 95 -250
rect 180 -280 195 -250
rect 80 -295 195 -280
<< nsubdiff >>
rect 70 375 220 385
rect 70 310 85 375
rect 205 310 220 375
rect 70 295 220 310
<< psubdiffcont >>
rect 95 -280 180 -250
<< nsubdiffcont >>
rect 85 310 205 375
<< poly >>
rect 130 205 145 260
rect 130 -30 145 -5
rect 65 -40 145 -30
rect 65 -70 75 -40
rect 105 -70 145 -40
rect 65 -80 145 -70
rect 200 -40 250 -30
rect 200 -70 210 -40
rect 240 -70 250 -40
rect 200 -80 250 -70
rect 130 -100 145 -80
rect 130 -215 145 -200
<< polycont >>
rect 75 -70 105 -40
rect 210 -70 240 -40
<< locali >>
rect 70 380 220 385
rect 70 375 100 380
rect 170 375 220 380
rect 70 310 85 375
rect 205 310 220 375
rect 70 300 100 310
rect 170 300 220 310
rect 70 295 220 300
rect 85 205 125 295
rect 80 195 125 205
rect 80 5 90 195
rect 115 5 125 195
rect 80 -5 125 5
rect 150 195 195 205
rect 150 5 160 195
rect 185 5 195 195
rect 150 -5 195 5
rect 155 -30 185 -5
rect 65 -40 115 -30
rect 65 -70 75 -40
rect 105 -70 115 -40
rect 65 -80 115 -70
rect 155 -40 250 -30
rect 155 -70 210 -40
rect 240 -70 250 -40
rect 155 -80 250 -70
rect 155 -100 185 -80
rect 85 -110 125 -100
rect 85 -190 95 -110
rect 115 -190 125 -110
rect 85 -200 125 -190
rect 150 -110 190 -100
rect 150 -190 160 -110
rect 180 -190 190 -110
rect 150 -200 190 -190
rect 90 -240 120 -200
rect 85 -250 115 -240
rect 160 -250 190 -240
rect 85 -280 95 -250
rect 180 -280 190 -250
rect 85 -285 115 -280
rect 160 -285 190 -280
rect 85 -290 190 -285
<< viali >>
rect 100 375 170 380
rect 100 310 170 375
rect 100 300 170 310
rect 75 -70 105 -40
rect 210 -70 240 -40
rect 115 -250 160 -240
rect 115 -280 160 -250
rect 115 -285 160 -280
<< metal1 >>
rect -240 380 545 385
rect -240 300 100 380
rect 170 300 545 380
rect -240 295 545 300
rect -210 -40 115 -30
rect -210 -70 75 -40
rect 105 -70 115 -40
rect -210 -80 115 -70
rect 155 -40 530 -30
rect 155 -70 210 -40
rect 240 -70 530 -40
rect 155 -80 530 -70
rect -220 -240 525 -235
rect -220 -285 115 -240
rect 160 -285 525 -240
rect -220 -295 525 -285
<< labels >>
rlabel metal1 450 325 450 325 1 vdd
rlabel metal1 500 -70 510 -45 1 out
rlabel metal1 -190 -70 -180 -45 1 in
<< end >>
