** sch_path: /mnt/c/Users/NITHIN P/Inverter_tb.sch
**.subckt Inverter_tb
x2 VDD Vin Vout GND CmosInverter
Vin Vin GND PULSE(0 1.8 0 0.1n 0.1n 10n 20n 10)
Vdd VDD GND 1.8
C2 Vout GND 0.1p m=1
**** begin user architecture code


.lib /home/nithinpuru/pdk/volare/sky130/versions/cd1748bb197f9b7af62a54507de6624e30363943/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran .02n 40n
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  /mnt/c/Users/NITHIN P/CmosInverter.sym # of pins=4
** sym_path: /mnt/c/Users/NITHIN P/CmosInverter.sym
** sch_path: /mnt/c/Users/NITHIN P/CmosInverter.sch
.subckt CmosInverter VDD Vin Vout VSS
*.ipin Vin
*.ipin VDD
*.ipin VSS
*.opin Vout
XM3 Vout Vin VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
